module lookup_table(
	input		clk,
	input		rst,
	input		[7:0]lut_in,
	output	[31:0]lut_out
    );

wire		clk,rst;
wire		[7:0]lut_in;
reg		[31:0]lut_out;


always @(posedge clk)
begin
	if (rst) begin
	lut_out =0;
	end else begin
	case (lut_in)
		8'b00000000: lut_out = 32'b00000000000000000000000000000000; //0
		8'b00000001: lut_out = 32'b00111111111111111111111111111001; //1
		8'b00000010: lut_out = 32'b00111111111111111111111111100010; //2
		8'b00000011: lut_out = 32'b00111111111111111111111110111011; //3
		8'b00000100: lut_out = 32'b00111111111111111111111110000101; //4
		8'b00000101: lut_out = 32'b00111111111111111111111100111111; //5
		8'b00000110: lut_out = 32'b00111111111111111111111011101010; //6
		8'b00000111: lut_out = 32'b00111111111111111111111010000101; //7
		8'b00001000: lut_out = 32'b00111111111111111111111000010001; //8
		8'b00001001: lut_out = 32'b00111111111111111111110110001101; //9
		8'b00001010: lut_out = 32'b00111111111111111111110011111010; //10
		8'b00001011: lut_out = 32'b00111111111111111111110001010111; //11
		8'b00001100: lut_out = 32'b00111111111111111111101110100101; //12
		8'b00001101: lut_out = 32'b00111111111111111111101011100100; //13
		8'b00001110: lut_out = 32'b00111111111111111111101000010010; //14
		8'b00001111: lut_out = 32'b00111111111111111111100100110010; //15
		8'b00010000: lut_out = 32'b00111111111111111111100001000010; //16
		8'b00010001: lut_out = 32'b00111111111111111111011101000010; //17
		8'b00010010: lut_out = 32'b00111111111111111111011000110011; //18
		8'b00010011: lut_out = 32'b00111111111111111111010100010100; //19
		8'b00010100: lut_out = 32'b00111111111111111111001111100110; //20
		8'b00010101: lut_out = 32'b00111111111111111111001010101001; //21
		8'b00010110: lut_out = 32'b00111111111111111111000101011100; //22
		8'b00010111: lut_out = 32'b00111111111111111110111111111111; //23
		8'b00011000: lut_out = 32'b00111111111111111110111010010011; //24
		8'b00011001: lut_out = 32'b00111111111111111110110100011000; //25
		8'b00011010: lut_out = 32'b00111111111111111110101110001101; //26
		8'b00011011: lut_out = 32'b00111111111111111110100111110010; //27
		8'b00011100: lut_out = 32'b00111111111111111110100001001000; //28
		8'b00011101: lut_out = 32'b00111111111111111110011010001111; //29
		8'b00011110: lut_out = 32'b00111111111111111110010011000110; //30
		8'b00011111: lut_out = 32'b00111111111111111110001011101101; //31
		8'b00100000: lut_out = 32'b00111111111111111110000100000101; //32
		8'b00100001: lut_out = 32'b00111111111111111101111100001110; //33
		8'b00100010: lut_out = 32'b00111111111111111101110100000111; //34
		8'b00100011: lut_out = 32'b00111111111111111101101011110000; //35
		8'b00100100: lut_out = 32'b00111111111111111101100011001010; //36
		8'b00100101: lut_out = 32'b00111111111111111101011010010101; //37
		8'b00100110: lut_out = 32'b00111111111111111101010001010000; //38
		8'b00100111: lut_out = 32'b00111111111111111101000111111100; //39
		8'b00101000: lut_out = 32'b00111111111111111100111110011000; //40
		8'b00101001: lut_out = 32'b00111111111111111100110100100100; //41
		8'b00101010: lut_out = 32'b00111111111111111100101010100010; //42
		8'b00101011: lut_out = 32'b00111111111111111100100000001111; //43
		8'b00101100: lut_out = 32'b00111111111111111100010101101101; //44
		8'b00101101: lut_out = 32'b00111111111111111100001010111100; //45
		8'b00101110: lut_out = 32'b00111111111111111011111111111011; //46
		8'b00101111: lut_out = 32'b00111111111111111011110100101011; //47
		8'b00110000: lut_out = 32'b00111111111111111011101001001011; //48
		8'b00110001: lut_out = 32'b00111111111111111011011101011100; //49
		8'b00110010: lut_out = 32'b00111111111111111011010001011101; //50
		8'b00110011: lut_out = 32'b00111111111111111011000101001111; //51
		8'b00110100: lut_out = 32'b00111111111111111010111000110001; //52
		8'b00110101: lut_out = 32'b00111111111111111010101100000100; //53
		8'b00110110: lut_out = 32'b00111111111111111010011111000111; //54
		8'b00110111: lut_out = 32'b00111111111111111010010001111011; //55
		8'b00111000: lut_out = 32'b00111111111111111010000100011111; //56
		8'b00111001: lut_out = 32'b00111111111111111001110110110100; //57
		8'b00111010: lut_out = 32'b00111111111111111001101000111001; //58
		8'b00111011: lut_out = 32'b00111111111111111001011010101111; //59
		8'b00111100: lut_out = 32'b00111111111111111001001100010101; //60
		8'b00111101: lut_out = 32'b00111111111111111000111101101100; //61
		8'b00111110: lut_out = 32'b00111111111111111000101110110011; //62
		8'b00111111: lut_out = 32'b00111111111111111000011111101011; //63
		8'b01000000: lut_out = 32'b00111111111111111000010000010011; //64
		8'b01000001: lut_out = 32'b00111111111111111000000000101100; //65
		8'b01000010: lut_out = 32'b00111111111111110111110000110101; //66
		8'b01000011: lut_out = 32'b00111111111111110111100000101111; //67
		8'b01000100: lut_out = 32'b00111111111111110111010000011010; //68
		8'b01000101: lut_out = 32'b00111111111111110110111111110101; //69
		8'b01000110: lut_out = 32'b00111111111111110110101111000000; //70
		8'b01000111: lut_out = 32'b00111111111111110110011101111100; //71
		8'b01001000: lut_out = 32'b00111111111111110110001100101000; //72
		8'b01001001: lut_out = 32'b00111111111111110101111011000101; //73
		8'b01001010: lut_out = 32'b00111111111111110101101001010011; //74
		8'b01001011: lut_out = 32'b00111111111111110101010111010001; //75
		8'b01001100: lut_out = 32'b00111111111111110101000100111111; //76
		8'b01001101: lut_out = 32'b00111111111111110100110010011110; //77
		8'b01001110: lut_out = 32'b00111111111111110100011111101101; //78
		8'b01001111: lut_out = 32'b00111111111111110100001100101101; //79
		8'b01010000: lut_out = 32'b00111111111111110011111001011110; //80
		8'b01010001: lut_out = 32'b00111111111111110011100101111111; //81
		8'b01010010: lut_out = 32'b00111111111111110011010010010000; //82
		8'b01010011: lut_out = 32'b00111111111111110010111110010010; //83
		8'b01010100: lut_out = 32'b00111111111111110010101010000101; //84
		8'b01010101: lut_out = 32'b00111111111111110010010101101000; //85
		8'b01010110: lut_out = 32'b00111111111111110010000000111011; //86
		8'b01010111: lut_out = 32'b00111111111111110001101011111111; //87
		8'b01011000: lut_out = 32'b00111111111111110001010110110100; //88
		8'b01011001: lut_out = 32'b00111111111111110001000001011001; //89
		8'b01011010: lut_out = 32'b00111111111111110000101011101111; //90
		8'b01011011: lut_out = 32'b00111111111111110000010101110101; //91
		8'b01011100: lut_out = 32'b00111111111111101111111111101011; //92
		8'b01011101: lut_out = 32'b00111111111111101111101001010010; //93
		8'b01011110: lut_out = 32'b00111111111111101111010010101010; //94
		8'b01011111: lut_out = 32'b00111111111111101110111011110010; //95
		8'b01100000: lut_out = 32'b00111111111111101110100100101011; //96
		8'b01100001: lut_out = 32'b00111111111111101110001101010100; //97
		8'b01100010: lut_out = 32'b00111111111111101101110101101110; //98
		8'b01100011: lut_out = 32'b00111111111111101101011101111000; //99
		8'b01100100: lut_out = 32'b00111111111111101101000101110010; //100
		8'b01100101: lut_out = 32'b00111111111111101100101101011110; //101
		8'b01100110: lut_out = 32'b00111111111111101100010100111001; //102
		8'b01100111: lut_out = 32'b00111111111111101011111100000101; //103
		8'b01101000: lut_out = 32'b00111111111111101011100011000010; //104
		8'b01101001: lut_out = 32'b00111111111111101011001001101111; //105
		8'b01101010: lut_out = 32'b00111111111111101010110000001101; //106
		8'b01101011: lut_out = 32'b00111111111111101010010110011011; //107
		8'b01101100: lut_out = 32'b00111111111111101001111100011010; //108
		8'b01101101: lut_out = 32'b00111111111111101001100010001001; //109
		8'b01101110: lut_out = 32'b00111111111111101001000111101001; //110
		8'b01101111: lut_out = 32'b00111111111111101000101100111001; //111
		8'b01110000: lut_out = 32'b00111111111111101000010001111010; //112
		8'b01110001: lut_out = 32'b00111111111111100111110110101011; //113
		8'b01110010: lut_out = 32'b00111111111111100111011011001101; //114
		8'b01110011: lut_out = 32'b00111111111111100110111111011111; //115
		8'b01110100: lut_out = 32'b00111111111111100110100011100010; //116
		8'b01110101: lut_out = 32'b00111111111111100110000111010110; //117
		8'b01110110: lut_out = 32'b00111111111111100101101010111001; //118
		8'b01110111: lut_out = 32'b00111111111111100101001110001110; //119
		8'b01111000: lut_out = 32'b00111111111111100100110001010011; //120
		8'b01111001: lut_out = 32'b00111111111111100100010100001000; //121
		8'b01111010: lut_out = 32'b00111111111111100011110110101110; //122
		8'b01111011: lut_out = 32'b00111111111111100011011001000100; //123
		8'b01111100: lut_out = 32'b00111111111111100010111011001011; //124
		8'b01111101: lut_out = 32'b00111111111111100010011101000010; //125
		8'b01111110: lut_out = 32'b00111111111111100001111110101010; //126
		8'b01111111: lut_out = 32'b00111111111111100001100000000011; //127
		8'b10000000: lut_out = 32'b00111111111111100001000001001100; //128
		8'b10000001: lut_out = 32'b00111111111111100000100010000101; //129
		8'b10000010: lut_out = 32'b00111111111111100000000010101111; //130
		8'b10000011: lut_out = 32'b00111111111111011111100011001010; //131
		8'b10000100: lut_out = 32'b00111111111111011111000011010100; //132
		8'b10000101: lut_out = 32'b00111111111111011110100011010000; //133
		8'b10000110: lut_out = 32'b00111111111111011110000010111100; //134
		8'b10000111: lut_out = 32'b00111111111111011101100010011000; //135
		8'b10001000: lut_out = 32'b00111111111111011101000001100101; //136
		8'b10001001: lut_out = 32'b00111111111111011100100000100011; //137
		8'b10001010: lut_out = 32'b00111111111111011011111111010001; //138
		8'b10001011: lut_out = 32'b00111111111111011011011101101111; //139
		8'b10001100: lut_out = 32'b00111111111111011010111011111110; //140
		8'b10001101: lut_out = 32'b00111111111111011010011001111110; //141
		8'b10001110: lut_out = 32'b00111111111111011001110111101110; //142
		8'b10001111: lut_out = 32'b00111111111111011001010101001111; //143
		8'b10010000: lut_out = 32'b00111111111111011000110010100000; //144
		8'b10010001: lut_out = 32'b00111111111111011000001111100001; //145
		8'b10010010: lut_out = 32'b00111111111111010111101100010011; //146
		8'b10010011: lut_out = 32'b00111111111111010111001000110110; //147
		8'b10010100: lut_out = 32'b00111111111111010110100101001001; //148
		8'b10010101: lut_out = 32'b00111111111111010110000001001101; //149
		8'b10010110: lut_out = 32'b00111111111111010101011101000001; //150
		8'b10010111: lut_out = 32'b00111111111111010100111000100101; //151
		8'b10011000: lut_out = 32'b00111111111111010100010011111011; //152
		8'b10011001: lut_out = 32'b00111111111111010011101111000000; //153
		8'b10011010: lut_out = 32'b00111111111111010011001001110110; //154
		8'b10011011: lut_out = 32'b00111111111111010010100100011101; //155
		8'b10011100: lut_out = 32'b00111111111111010001111110110100; //156
		8'b10011101: lut_out = 32'b00111111111111010001011000111100; //157
		8'b10011110: lut_out = 32'b00111111111111010000110010110100; //158
		8'b10011111: lut_out = 32'b00111111111111010000001100011101; //159
		8'b10100000: lut_out = 32'b00111111111111001111100101110110; //160
		8'b10100001: lut_out = 32'b00111111111111001110111111000000; //161
		8'b10100010: lut_out = 32'b00111111111111001110010111111010; //162
		8'b10100011: lut_out = 32'b00111111111111001101110000100101; //163
		8'b10100100: lut_out = 32'b00111111111111001101001001000000; //164
		8'b10100101: lut_out = 32'b00111111111111001100100001001100; //165
		8'b10100110: lut_out = 32'b00111111111111001011111001001000; //166
		8'b10100111: lut_out = 32'b00111111111111001011010000110101; //167
		8'b10101000: lut_out = 32'b00111111111111001010101000010010; //168
		8'b10101001: lut_out = 32'b00111111111111001001111111100000; //169
		8'b10101010: lut_out = 32'b00111111111111001001010110011110; //170
		8'b10101011: lut_out = 32'b00111111111111001000101101001101; //171
		8'b10101100: lut_out = 32'b00111111111111001000000011101100; //172
		8'b10101101: lut_out = 32'b00111111111111000111011001111100; //173
		8'b10101110: lut_out = 32'b00111111111111000110101111111100; //174
		8'b10101111: lut_out = 32'b00111111111111000110000101101101; //175
		8'b10110000: lut_out = 32'b00111111111111000101011011001111; //176
		8'b10110001: lut_out = 32'b00111111111111000100110000100001; //177
		8'b10110010: lut_out = 32'b00111111111111000100000101100011; //178
		8'b10110011: lut_out = 32'b00111111111111000011011010010110; //179
		8'b10110100: lut_out = 32'b00111111111111000010101110111001; //180
		8'b10110101: lut_out = 32'b00111111111111000010000011001101; //181
		8'b10110110: lut_out = 32'b00111111111111000001010111010010; //182
		8'b10110111: lut_out = 32'b00111111111111000000101011000110; //183
		8'b10111000: lut_out = 32'b00111111111110111111111110101100; //184
		8'b10111001: lut_out = 32'b00111111111110111111010010000010; //185
		8'b10111010: lut_out = 32'b00111111111110111110100101001000; //186
		8'b10111011: lut_out = 32'b00111111111110111101110111111111; //187
		8'b10111100: lut_out = 32'b00111111111110111101001010100111; //188
		8'b10111101: lut_out = 32'b00111111111110111100011100111111; //189
		8'b10111110: lut_out = 32'b00111111111110111011101111000111; //190
		8'b10111111: lut_out = 32'b00111111111110111011000001000000; //191
		8'b11000000: lut_out = 32'b00111111111110111010010010101010; //192
		8'b11000001: lut_out = 32'b00111111111110111001100100000100; //193
		8'b11000010: lut_out = 32'b00111111111110111000110101001110; //194
		8'b11000011: lut_out = 32'b00111111111110111000000110001001; //195
		8'b11000100: lut_out = 32'b00111111111110110111010110110101; //196
		8'b11000101: lut_out = 32'b00111111111110110110100111010001; //197
		8'b11000110: lut_out = 32'b00111111111110110101110111011101; //198
		8'b11000111: lut_out = 32'b00111111111110110101000111011011; //199
		8'b11001000: lut_out = 32'b00111111111110110100010111001000; //200
		8'b11001001: lut_out = 32'b00111111111110110011100110100110; //201
		8'b11001010: lut_out = 32'b00111111111110110010110101110101; //202
		8'b11001011: lut_out = 32'b00111111111110110010000100110100; //203
		8'b11001100: lut_out = 32'b00111111111110110001010011100100; //204
		8'b11001101: lut_out = 32'b00111111111110110000100010000100; //205
		8'b11001110: lut_out = 32'b00111111111110101111110000010100; //206
		8'b11001111: lut_out = 32'b00111111111110101110111110010101; //207
		8'b11010000: lut_out = 32'b00111111111110101110001100000111; //208
		8'b11010001: lut_out = 32'b00111111111110101101011001101001; //209
		8'b11010010: lut_out = 32'b00111111111110101100100110111100; //210
		8'b11010011: lut_out = 32'b00111111111110101011110011111111; //211
		8'b11010100: lut_out = 32'b00111111111110101011000000110011; //212
		8'b11010101: lut_out = 32'b00111111111110101010001101010111; //213
		8'b11010110: lut_out = 32'b00111111111110101001011001101100; //214
		8'b11010111: lut_out = 32'b00111111111110101000100101110001; //215
		8'b11011000: lut_out = 32'b00111111111110100111110001100111; //216
		8'b11011001: lut_out = 32'b00111111111110100110111101001101; //217
		8'b11011010: lut_out = 32'b00111111111110100110001000100100; //218
		8'b11011011: lut_out = 32'b00111111111110100101010011101011; //219
		8'b11011100: lut_out = 32'b00111111111110100100011110100011; //220
		8'b11011101: lut_out = 32'b00111111111110100011101001001011; //221
		8'b11011110: lut_out = 32'b00111111111110100010110011100100; //222
		8'b11011111: lut_out = 32'b00111111111110100001111101101101; //223
		8'b11100000: lut_out = 32'b00111111111110100001000111100111; //224
		8'b11100001: lut_out = 32'b00111111111110100000010001010001; //225
		8'b11100010: lut_out = 32'b00111111111110011111011010101100; //226
		8'b11100011: lut_out = 32'b00111111111110011110100011110111; //227
		8'b11100100: lut_out = 32'b00111111111110011101101100110011; //228
		8'b11100101: lut_out = 32'b00111111111110011100110101011111; //229
		8'b11100110: lut_out = 32'b00111111111110011011111101111100; //230
		8'b11100111: lut_out = 32'b00111111111110011011000110001010; //231
		8'b11101000: lut_out = 32'b00111111111110011010001110001000; //232
		8'b11101001: lut_out = 32'b00111111111110011001010101110110; //233
		8'b11101010: lut_out = 32'b00111111111110011000011101010101; //234
		8'b11101011: lut_out = 32'b00111111111110010111100100100100; //235
		8'b11101100: lut_out = 32'b00111111111110010110101011100100; //236
		8'b11101101: lut_out = 32'b00111111111110010101110010010101; //237
		8'b11101110: lut_out = 32'b00111111111110010100111000110101; //238
		8'b11101111: lut_out = 32'b00111111111110010011111111000111; //239
		8'b11110000: lut_out = 32'b00111111111110010011000101001001; //240
		8'b11110001: lut_out = 32'b00111111111110010010001010111011; //241
		8'b11110010: lut_out = 32'b00111111111110010001010000011110; //242
		8'b11110011: lut_out = 32'b00111111111110010000010101110010; //243
		8'b11110100: lut_out = 32'b00111111111110001111011010110110; //244
		8'b11110101: lut_out = 32'b00111111111110001110011111101010; //245
		8'b11110110: lut_out = 32'b00111111111110001101100100001111; //246
		8'b11110111: lut_out = 32'b00111111111110001100101000100101; //247
		8'b11111000: lut_out = 32'b00111111111110001011101100101011; //248
		8'b11111001: lut_out = 32'b00111111111110001010110000100001; //249
		8'b11111010: lut_out = 32'b00111111111110001001110100001000; //250
		8'b11111011: lut_out = 32'b00111111111110001000110111100000; //251
		8'b11111100: lut_out = 32'b00111111111110000111111010101000; //252
		8'b11111101: lut_out = 32'b00111111111110000110111101100001; //253
		8'b11111110: lut_out = 32'b00111111111110000110000000001010; //254
		8'b11111111: lut_out = 32'b00111111111110000101000010100011; //255
		default	  : lut_out = 32'b00000000000000000000000000000000;	
	endcase
	end
end


endmodule
